#must fail
