../microwatt/insn_helpers.vhdl