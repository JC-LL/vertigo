../microwatt/wishbone_arbiter.vhdl