../microwatt/logical.vhdl