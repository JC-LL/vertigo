../microwatt/sim_console.vhdl