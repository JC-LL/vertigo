package body lfsr_pkg is

    function func (x:boolean) return boolean is
    begin
        
        v11 := a;
	
    end function;

    
end package body;


    
