
architecture rtl of aggregate_2 is

begin
  bus_data_a2p <= x"0000000" & "000" & ifregs.ctrl;
end rtl;
