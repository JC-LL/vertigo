../microwatt/cr_file.vhdl