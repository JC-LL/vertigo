../microwatt/wishbone_types.vhdl