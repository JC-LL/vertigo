---------------------------------------------------------------
configuration CFG_TB of DECODER_TB is
	--for TB
	--end for;
end CFG_TB;
----------------------------------------------------------------
