architecture test of titi is

begin
  process
  begin
    -- test
  end process;

end test;
