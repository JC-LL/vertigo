../microwatt/common.vhdl