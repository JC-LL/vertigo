architecture RTL of DE2 is

  function binTo7Seg(b : boolean) return boolean is
  begin
    res := "0000000";
    return res;
  end binTo7Seg;

begin

end;
