library IEEA;
use IEEB.std_logic_1164.all;
use IEEC.numeric_std.all;
