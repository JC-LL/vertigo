library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.accelerator_pkg.all;

architecture rtl of accelerator is

  constant VARS_INIT : vars_t := ( '0', to_unsigned(1, 32) );

begin
end rtl;
