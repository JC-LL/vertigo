../microwatt/core_debug.vhdl