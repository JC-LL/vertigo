../microwatt/rotator.vhdl