library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.accelerator_pkg.all;

architecture rtl of accelerator is
  signal s : unsigned := to_unsigned(0, 32);
begin
end rtl;
