../microwatt/plru_tb.vhdl