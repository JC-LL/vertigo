../microwatt/cr_hazard.vhdl