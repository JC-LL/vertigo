f(x,y)
