( a => '0', to_unsigned(1, 32) )
