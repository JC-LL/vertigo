../microwatt/glibc_random_helpers.vhdl