
architecture test of aggregate_2 is

begin
  test.a.b.c <= '0';
end rtl;
