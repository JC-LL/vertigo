../microwatt/icache_tb.vhdl