( '0', "0000", x"FFFF", 42)
