entity test is
end;

architecture test_var of test is

  type TestIt is array(natural range <>) of boolean;

begin
end test_var;
