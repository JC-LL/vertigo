package lfsr_pkg is

 function test(a,b: boolean;
               c : integer;
               d : std_logic_vector(1 downto 0)) return boolean;
    
end package;


    
