../microwatt/gpr_hazard.vhdl