../microwatt/decode2.vhdl