../microwatt/utils.vhdl