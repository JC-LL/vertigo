
architecture test_var of test is
  
  type mem2 is array(1 to 100) of integer;

begin
end test_var;

