
package ALU_package is

	procedure check(a : integer);
    
end ALU_package;  

