../microwatt/divider.vhdl