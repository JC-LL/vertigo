
architecture test_var of test is
  
  type mem2 is array(1 to 100) of integer;

begin  -- test_var
  
  test : process
    --type mem2 is array(1 to 100) of integer;
    --type TestIt is array(natural range <>) of boolean;
    --type    Mem is array (natural range <>, natural range <>) of integer;
  begin  
  end process test;
  
end test_var;

