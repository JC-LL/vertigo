package body lfsr_pkg is

 function t(a: boolean) return boolean is
   variable v1 : boolean;
 begin
   null; 
 end;
    
end package body;


    
