../microwatt/control.vhdl