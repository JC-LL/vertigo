../microwatt/dmi_dtm_tb.vhdl