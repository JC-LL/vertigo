../microwatt/wishbone_debug_master.vhdl