../microwatt/dmi_dtm_xilinx.vhdl