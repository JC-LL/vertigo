../microwatt/sim_uart.vhdl