../microwatt/core_tb.vhdl