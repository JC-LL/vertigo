../microwatt/sim_bram_helpers.vhdl