../microwatt/fetch2.vhdl