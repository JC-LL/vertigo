../microwatt/rotator_tb.vhdl