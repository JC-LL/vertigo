../microwatt/countzero.vhdl