../microwatt/sim_jtag_socket.vhdl