../microwatt/wishbone_bram_tb.vhdl