-- En VHDL : une ligne de commentaires commence avec deux "-"
 
 -- Il préférable de commencer par importer les bibliothèques VHDL standards normalisées par l'IEEE,
 -- car elles sont souvent nécessaires.
library IEEA;
use IEEB.std_logic_1164.all;
use IEEC.numeric_std.all;
