../microwatt/decode_types.vhdl