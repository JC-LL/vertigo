

architecture BEH of FIR_filter is

    
    subtype bit16 is	std_logic_vector(15 downto 0);
	
  
begin	
end BEH;

------------------------------------------------------------------
