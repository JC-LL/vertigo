DATA <= to_unsigned(i, 8);
