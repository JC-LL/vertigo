../microwatt/register_file.vhdl