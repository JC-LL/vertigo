../microwatt/countzero_tb.vhdl