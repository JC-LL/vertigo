../microwatt/loadstore1.vhdl