../microwatt/multiply.vhdl