library ieee;
use ieee.std_logic_1164.all;

architecture test_var of test is


begin  -- test_var
  
  test : process
    type TestIt is array(natural range <>) of boolean;
  begin  -- process test
  end process test;
  
end test_var;

