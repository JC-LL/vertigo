../microwatt/fetch1.vhdl