../microwatt/sim_jtag.vhdl