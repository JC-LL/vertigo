../microwatt/sim_bram.vhdl