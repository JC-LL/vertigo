../microwatt/divider_tb.vhdl