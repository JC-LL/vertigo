../microwatt/crhelpers.vhdl