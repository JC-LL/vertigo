../microwatt/glibc_random.vhdl