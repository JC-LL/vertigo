../microwatt/dcache.vhdl