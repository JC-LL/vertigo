../microwatt/writeback.vhdl