../microwatt/wishbone_bram_wrapper.vhdl