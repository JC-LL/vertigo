../microwatt/ppc_fx_insns.vhdl