 entity logique_4_vers_1 is 
 end logique_4_vers_1;
