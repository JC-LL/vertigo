../microwatt/execute1.vhdl