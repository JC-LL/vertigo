

package body test is

    function f (a, b :integer) return boolean is
    begin
      return true;
    end function;

end package body;


    
