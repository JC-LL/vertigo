../microwatt/helpers.vhdl