-- Première architecture concurrente décrivant un mux :
 ARCHITECTURE mux_4_vers_1 OF logique_4_vers_1 IS
 
 BEGIN

 END mux_4_vers_1;
