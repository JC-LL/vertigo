../microwatt/decode1.vhdl