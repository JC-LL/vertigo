../microwatt/icache.vhdl