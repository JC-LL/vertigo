../microwatt/cache_ram.vhdl