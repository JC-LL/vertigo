../microwatt/dmi_dtm_dummy.vhdl