../microwatt/multiply_tb.vhdl