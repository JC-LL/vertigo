../microwatt/plru.vhdl