( a => '0')
