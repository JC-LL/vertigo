

architecture BEH of FIR_filter is  
begin	
end BEH;

--------------