Output_X(i) <= Input_X(i+8) after 5 ns;
