
architecture test_var of test is
  
begin  
  
  test : process
  begin  
  end process test;
  
end test_var;

