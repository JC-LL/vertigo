../microwatt/core.vhdl