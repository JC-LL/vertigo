../microwatt/dcache_tb.vhdl