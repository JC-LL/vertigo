../microwatt/soc.vhdl